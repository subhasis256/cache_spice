.param Wn=16.50
.param Wp=49.50
.param Wload=176.467
.param Rload=3.584
.include "inv.ckt"
