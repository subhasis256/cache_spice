.param Wn=224.14
.param Wp=672.41
.param Wload=2823.478
.param Rload=57.344
.include "inv.ckt"
