.param Wn=83.26
.param Wp=249.79
.param Wload=705.869
.param Rload=14.336
.include "inv.ckt"
