.param Wn=21.18
.param Wp=63.54
.param Wload=176.467
.param Rload=3.584
.include "inv.ckt"
