.param Nw=1024
.param Nh=256
