.param Nw=128
.param Nh=16
