.param Nw=16
.param Nh=16
