.param Nw=256
.param Nh=256
