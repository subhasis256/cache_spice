.param Wn=97.48
.param Wp=292.44
.param Wload=705.869
.param Rload=14.336
.include "inv.ckt"
