.param Rperl=4000k
.param Lperl=1.952u
.param Cperl=297.5p
.param length=171.1u
.param iscale=200

